module cmp

pub enum Ordering {
	less
	equal
	greater
}